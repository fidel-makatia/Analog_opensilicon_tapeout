* ============================================================================
* OTA AC Gain/Phase Analysis Testbench
* ============================================================================
* Measures open-loop gain, unity-gain bandwidth, and phase margin
*
* Usage: ngspice -b ota_tb_ac.spice
* ============================================================================

.lib $PDK_ROOT/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.include "ota.spice"

* ---- Power Supply ----
VDD VDD 0 1.8
VSS VSS 0 0

* ---- Bias with AC stimulus on VIN+ ----
VINP VINP 0 DC 0.9 AC 1
VINN VINN 0 0.9

* ---- External reference current (10uA from VDD into IREF node) ----
IIREF VDD IREF 10u

* ---- Load capacitor ----
CL VOUT VSS 1p

* ---- Instantiate OTA ----
XOTA VINP VINN VOUT VDD VSS IREF ota

* ---- AC Analysis: 100 points/decade, 1Hz to 1GHz ----
.ac dec 100 1 1G

.control
  run
  echo ""
  echo "============================================================"
  echo "  OTA AC Analysis Results"
  echo "============================================================"

  * Measure DC gain
  meas ac dc_gain find vdb(VOUT) at=10
  echo ""

  * Measure unity-gain bandwidth
  meas ac ugb when vdb(VOUT)=0
  echo ""

  * Measure phase margin at UGB
  meas ac phase_at_ugb find vp(VOUT) when vdb(VOUT)=0
  echo ""

  echo "  Target: DC Gain 20-35 dB, UGB 1-3 MHz"
  echo "============================================================"

  * Save Bode data
  wrdata ../outputs/ac_bode.csv vdb(VOUT) vp(VOUT)
  echo "  Bode data saved to outputs/ac_bode.csv"
  quit
.endc

.end
